<svg xmlns="http://www.w3.org/2000/svg" width="480" height="351" class="">
    <defs>
        <style/>
    </defs>
    <style>@keyframes animation-gauge{0%{stroke-dasharray:0 329}}@keyframes animation-fade{0%{opacity:0}to{opacity:1}}@keyframes animation-rainbow{0%,to{color:#7f00ff;fill:#7f00ff}14%{color:#a933ff;fill:#a933ff}29%{color:#007fff;fill:#007fff}43%{color:#00ff7f;fill:#00ff7f}57%{color:#ff0;fill:#ff0}71%{color:#ff7f00;fill:#ff7f00}86%{color:red;fill:red}}svg{font-family:-apple-system,BlinkMacSystemFont,Segoe UI,Helvetica,Arial,sans-serif,Apple Color Emoji,Segoe UI Emoji;color:#777}h2,h3{margin:8px 0 2px;padding:0;color:#0366d6;font-weight:400}h2 svg,h3 svg{fill:currentColor}h2{font-size:16px}h3,svg{font-size:14px}section&gt;.field{margin-left:5px;margin-right:5px}.field{display:flex;align-items:center;margin-bottom:2px;white-space:nowrap}.field svg{margin:0 8px;fill:#959da5;flex-shrink:0}.row{display:flex;flex-wrap:wrap}.row section{flex:1 1 0}.column{display:flex;flex-direction:column;align-items:center}#metrics-end,.fill-width{width:100%}.calendar.field{margin:4px 0 4px 7px}.calendar .day{outline:1px solid rgba(27,31,35,.04);outline-offset:-1px}svg.bar{margin:4px 0}.field.language{margin:0 8px;flex-grow:0}.field.language.details,.field.language.details small{display:flex;justify-content:space-between}.field.language.details small{color:#666;text-align:right}.field.language.details small&gt;*,.field.language.details&gt;*{flex:1 1 0}.field.language.details small&gt;:not(:last-child){margin-right:6px}.footnote{width:100%;justify-content:flex-end;font-size:12px}.chartist .ct-post{fill:rgba(127,127,127,.8)!important;color:rgba(127,127,127,.8)!important;font-size:9px;text-anchor:middle}:root{--color-calendar-graph-day-bg:#ebedf0;--color-calendar-graph-day-border:rgba(27,31,35,0.06);--color-calendar-graph-day-L1-bg:#9be9a8;--color-calendar-graph-day-L2-bg:#40c463;--color-calendar-graph-day-L3-bg:#30a14e;--color-calendar-graph-day-L4-bg:#216e39;--color-calendar-halloween-graph-day-L1-bg:#ffee4a;--color-calendar-halloween-graph-day-L2-bg:#ffc501;--color-calendar-halloween-graph-day-L3-bg:#fe9600;--color-calendar-halloween-graph-day-L4-bg:#03001c;--color-calendar-graph-day-L4-border:rgba(27,31,35,0.06);--color-calendar-graph-day-L3-border:rgba(27,31,35,0.06);--color-calendar-graph-day-L2-border:rgba(27,31,35,0.06);--color-calendar-graph-day-L1-border:rgba(27,31,35,0.06)}</style>
    <style/>
    <foreignObject x="0" y="0" width="100%" height="100%">
        <div xmlns="http://www.w3.org/1999/xhtml" xmlns:xlink="http://www.w3.org/1999/xlink" class="items-wrapper">
            <section>
                <h2 class="field">
                    <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                        <path fill-rule="evenodd" d="M1.5 2.75a.25.25 0 01.25-.25h12.5a.25.25 0 01.25.25v8.5a.25.25 0 01-.25.25h-6.5a.75.75 0 00-.53.22L4.5 14.44v-2.19a.75.75 0 00-.75-.75h-2a.25.25 0 01-.25-.25v-8.5zM1.75 1A1.75 1.75 0 000 2.75v8.5C0 12.216.784 13 1.75 13H3v1.543a1.457 1.457 0 002.487 1.03L8.061 13h6.189A1.75 1.75 0 0016 11.25v-8.5A1.75 1.75 0 0014.25 1H1.75zm5.03 3.47a.75.75 0 010 1.06L5.31 7l1.47 1.47a.75.75 0 01-1.06 1.06l-2-2a.75.75 0 010-1.06l2-2a.75.75 0 011.06 0zm2.44 0a.75.75 0 000 1.06L10.69 7 9.22 8.47a.75.75 0 001.06 1.06l2-2a.75.75 0 000-1.06l-2-2a.75.75 0 00-1.06 0z"/>
                    </svg>
                    2 Languages
                </h2>
            </section>
            <section class="column">
                <h3 class="field">Most used languages</h3>
                <small>estimation from 24 edited files from 50 commits</small>
                <svg class="bar" xmlns="http://www.w3.org/2000/svg" width="460" height="8">
                    <mask id="languages-bar">
                        <rect x="0" y="0" width="460" height="8" fill="white" rx="5"/>
                    </mask>
                    <rect mask="url(#languages-bar)" x="0" y="0" width="0" height="8" fill="#d1d5da"/>
                    <rect mask="url(#languages-bar)" x="0" y="0" width="460" height="8" fill="#f1e05a"/>
                </svg>
                <div class="row fill-width">
                    <section>
                        <div class="field language details">
                            <div class="field">
                                <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                    <path fill="#f1e05a" fill-rule="evenodd" d="M8 4a4 4 0 100 8 4 4 0 000-8z"/>
                                </svg>
                                JavaScript
                            </div>
                            <small>
                                <div>476 lines</div>
                                <div>11.8 kB</div>
                            </small>
                        </div>
                    </section>
                    <section>
                    </section>
                </div>
                <div class="row footnote">
                    <div class="field">
                        <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                            <path fill-rule="evenodd" d="M9.585.52a2.678 2.678 0 00-3.17 0l-.928.68a1.178 1.178 0 01-.518.215L3.83 1.59a2.678 2.678 0 00-2.24 2.24l-.175 1.14a1.178 1.178 0 01-.215.518l-.68.928a2.678 2.678 0 000 3.17l.68.928c.113.153.186.33.215.518l.175 1.138a2.678 2.678 0 002.24 2.24l1.138.175c.187.029.365.102.518.215l.928.68a2.678 2.678 0 003.17 0l.928-.68a1.17 1.17 0 01.518-.215l1.138-.175a2.678 2.678 0 002.241-2.241l.175-1.138c.029-.187.102-.365.215-.518l.68-.928a2.678 2.678 0 000-3.17l-.68-.928a1.179 1.179 0 01-.215-.518L14.41 3.83a2.678 2.678 0 00-2.24-2.24l-1.138-.175a1.179 1.179 0 01-.518-.215L9.585.52zM7.303 1.728c.415-.305.98-.305 1.394 0l.928.68c.348.256.752.423 1.18.489l1.136.174c.51.078.909.478.987.987l.174 1.137c.066.427.233.831.489 1.18l.68.927c.305.415.305.98 0 1.394l-.68.928a2.678 2.678 0 00-.489 1.18l-.174 1.136a1.178 1.178 0 01-.987.987l-1.137.174a2.678 2.678 0 00-1.18.489l-.927.68c-.415.305-.98.305-1.394 0l-.928-.68a2.678 2.678 0 00-1.18-.489l-1.136-.174a1.178 1.178 0 01-.987-.987l-.174-1.137a2.678 2.678 0 00-.489-1.18l-.68-.927a1.178 1.178 0 010-1.394l.68-.928c.256-.348.423-.752.489-1.18l.174-1.136c.078-.51.478-.909.987-.987l1.137-.174a2.678 2.678 0 001.18-.489l.927-.68zM11.28 6.78a.75.75 0 00-1.06-1.06L7 8.94 5.78 7.72a.75.75 0 00-1.06 1.06l1.75 1.75a.75.75 0 001.06 0l3.75-3.75z"/>
                        </svg>
                        48 commits verified by GPG
                    </div>
                </div>
            </section>
            <section>
                <h2 class="field">
                    <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                        <path fill-rule="evenodd" d="M4.75 0a.75.75 0 01.75.75V2h5V.75a.75.75 0 011.5 0V2h1.25c.966 0 1.75.784 1.75 1.75v10.5A1.75 1.75 0 0113.25 16H2.75A1.75 1.75 0 011 14.25V3.75C1 2.784 1.784 2 2.75 2H4V.75A.75.75 0 014.75 0zm0 3.5h8.5a.25.25 0 01.25.25V6h-11V3.75a.25.25 0 01.25-.25h2zm-2.25 4v6.75c0 .138.112.25.25.25h10.5a.25.25 0 00.25-.25V7.5h-11z"/>
                    </svg>
                    Contributions calendar
                </h2>
                <div class="row">
                    <section>
                    </section>
                    <section>
                        <h3 class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path fill-rule="evenodd" d="M7.75 14A1.75 1.75 0 016 12.25v-8.5C6 2.784 6.784 2 7.75 2h6.5c.966 0 1.75.784 1.75 1.75v8.5A1.75 1.75 0 0114.25 14h-6.5zm-.25-1.75c0 .138.112.25.25.25h6.5a.25.25 0 00.25-.25v-8.5a.25.25 0 00-.25-.25h-6.5a.25.25 0 00-.25.25v8.5zM4.9 3.508a.75.75 0 01-.274 1.025.25.25 0 00-.126.217v6.5a.25.25 0 00.126.217.75.75 0 01-.752 1.298A1.75 1.75 0 013 11.25v-6.5c0-.649.353-1.214.874-1.516a.75.75 0 011.025.274zM1.625 5.533a.75.75 0 10-.752-1.299A1.75 1.75 0 000 5.75v4.5c0 .649.353 1.214.874 1.515a.75.75 0 10.752-1.298.25.25 0 01-.126-.217v-4.5a.25.25 0 01.126-.217z"/>
                            </svg>
                            Commits streaks
                        </h3>
                        <div class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path fill-rule="evenodd" d="M7.998 14.5c2.832 0 5-1.98 5-4.5 0-1.463-.68-2.19-1.879-3.383l-.036-.037c-1.013-1.008-2.3-2.29-2.834-4.434-.322.256-.63.579-.864.953-.432.696-.621 1.58-.046 2.73.473.947.67 2.284-.278 3.232-.61.61-1.545.84-2.403.633a2.788 2.788 0 01-1.436-.874A3.21 3.21 0 003 10c0 2.53 2.164 4.5 4.998 4.5zM9.533.753C9.496.34 9.16.009 8.77.146 7.035.75 4.34 3.187 5.997 6.5c.344.689.285 1.218.003 1.5-.419.419-1.54.487-2.04-.832-.173-.454-.659-.762-1.035-.454C2.036 7.44 1.5 8.702 1.5 10c0 3.512 2.998 6 6.498 6s6.5-2.5 6.5-6c0-2.137-1.128-3.26-2.312-4.438-1.19-1.184-2.436-2.425-2.653-4.81z"/>
                            </svg>
                            Current streak 1 day
                        </div>
                        <div class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path d="M8.5.75a.75.75 0 00-1.5 0v5.19L4.391 3.33a.75.75 0 10-1.06 1.061L5.939 7H.75a.75.75 0 000 1.5h5.19l-2.61 2.609a.75.75 0 101.061 1.06L7 9.561v5.189a.75.75 0 001.5 0V9.56l2.609 2.61a.75.75 0 101.06-1.061L9.561 8.5h5.189a.75.75 0 000-1.5H9.56l2.61-2.609a.75.75 0 00-1.061-1.06L8.5 5.939V.75z"/>
                            </svg>
                            Best streak 3 days
                        </div>
                        <h3 class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path fill-rule="evenodd" d="M10.5 7.75a2.5 2.5 0 11-5 0 2.5 2.5 0 015 0zm1.43.75a4.002 4.002 0 01-7.86 0H.75a.75.75 0 110-1.5h3.32a4.001 4.001 0 017.86 0h3.32a.75.75 0 110 1.5h-3.32z"/>
                            </svg>
                            Commits per day
                        </h3>
                        <div class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path d="M7.823 1.677L4.927 4.573A.25.25 0 005.104 5H7.25v3.236a.75.75 0 101.5 0V5h2.146a.25.25 0 00.177-.427L8.177 1.677a.25.25 0 00-.354 0zM13.75 11a.75.75 0 000 1.5h.5a.75.75 0 000-1.5h-.5zm-3.75.75a.75.75 0 01.75-.75h.5a.75.75 0 010 1.5h-.5a.75.75 0 01-.75-.75zM7.75 11a.75.75 0 000 1.5h.5a.75.75 0 000-1.5h-.5zM4 11.75a.75.75 0 01.75-.75h.5a.75.75 0 010 1.5h-.5a.75.75 0 01-.75-.75zM1.75 11a.75.75 0 000 1.5h.5a.75.75 0 000-1.5h-.5z"/>
                            </svg>
                            Highest in a day at 10
                        </div>
                        <div class="field">
                            <svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 16 16" width="16" height="16">
                                <path d="M10.896 2H8.75V.75a.75.75 0 00-1.5 0V2H5.104a.25.25 0 00-.177.427l2.896 2.896a.25.25 0 00.354 0l2.896-2.896A.25.25 0 0010.896 2zM8.75 15.25a.75.75 0 01-1.5 0V14H5.104a.25.25 0 01-.177-.427l2.896-2.896a.25.25 0 01.354 0l2.896 2.896a.25.25 0 01-.177.427H8.75v1.25zm-6.5-6.5a.75.75 0 000-1.5h-.5a.75.75 0 000 1.5h.5zM6 8a.75.75 0 01-.75.75h-.5a.75.75 0 010-1.5h.5A.75.75 0 016 8zm2.25.75a.75.75 0 000-1.5h-.5a.75.75 0 000 1.5h.5zM12 8a.75.75 0 01-.75.75h-.5a.75.75 0 010-1.5h.5A.75.75 0 0112 8zm2.25.75a.75.75 0 000-1.5h-.5a.75.75 0 000 1.5h.5z"/>
                            </svg>
                            Average per day at ~0.18
                        </div>
                    </section>
                </div>
                <svg version="1.1" xmlns="http://www.w3.org/2000/svg" style="margin-top: -130px;" viewBox="0,0 480,170">
                    <filter id="brightness1">
                        <feComponentTransfer>
                            <feFuncR type="linear" slope="0.6"/>
                            <feFuncG type="linear" slope="0.6"/>
                            <feFuncB type="linear" slope="0.6"/>
                        </feComponentTransfer>
                    </filter>
                    <filter id="brightness2">
                        <feComponentTransfer>
                            <feFuncR type="linear" slope="0.19999999999999996"/>
                            <feFuncG type="linear" slope="0.19999999999999996"/>
                            <feFuncB type="linear" slope="0.19999999999999996"/>
                        </feComponentTransfer>
                    </filter>
                    <g transform="scale(4) translate(12, 0)">
                        <g transform="translate(0, 0)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(1.7, 1)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(3.4, 2)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(5.1, 3)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(6.8, 4)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(8.5, 5)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(10.2, 6)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(11.9, 7)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(13.6, 8)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(15.299999999999999, 9)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.4)">
                                <path fill="#9be9a8" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#9be9a8" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6 0,1.6 z"/>
                                <path fill="#9be9a8" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.6 1.7,2.6 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 9)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,5 0,4 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,4 1.7,5 z"/>
                            </g>
                        </g>
                        <g transform="translate(17, 10)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(18.7, 11)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 8)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,5 0,4 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,4 1.7,5 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(20.4, 12)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(22.099999999999998, 13)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(23.8, 14)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(25.5, 15)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(27.2, 16)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(28.9, 17)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(30.599999999999998, 18)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 6)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,8 0,7 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,7 1.7,8 z"/>
                            </g>
                        </g>
                        <g transform="translate(32.3, 19)">
                            <g transform="translate(0, 5.4)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6 0,1.6 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.6 1.7,2.6 z"/>
                            </g>
                            <g transform="translate(-1.7, 5.800000000000001)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.2 0,2.2 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.2 1.7,3.2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(34, 20)">
                            <g transform="translate(0, 5.4)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6 0,1.6 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.6 1.7,2.6 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(35.699999999999996, 21)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 9.8)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.2 0,2.2 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.2 1.7,3.2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(37.4, 22)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(39.1, 23)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 8.4)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6 0,1.6 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.6 1.7,2.6 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(40.8, 24)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 7)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 9.4)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6 0,1.6 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.6 1.7,2.6 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 12)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                        </g>
                        <g transform="translate(42.5, 25)">
                            <g transform="translate(0, 6)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-1.7, 6.4)">
                                <path fill="#40c463" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#40c463" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2.6 0,1.6 z"/>
                                <path fill="#40c463" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1.6 1.7,2.6 z"/>
                            </g>
                            <g transform="translate(-3.4, 8)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-5.1, 9)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-6.8, 10)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-8.5, 11)">
                                <path fill="#ebedf0" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,2 0,1 z"/>
                                <path fill="#ebedf0" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,1 1.7,2 z"/>
                            </g>
                            <g transform="translate(-10.2, 10.2)">
                                <path fill="#216e39" d="M1.7,2 0,1 1.7,0 3.4,1 z"/>
                                <path fill="#216e39" filter="url(#brightness1)" d="M0,1 1.7,2 1.7,3.8 0,2.8 z"/>
                                <path fill="#216e39" filter="url(#brightness2)" d="M1.7,2 3.4,1 3.4,2.8 1.7,3.8 z"/>
                            </g>
                        </g>
                    </g>
                </svg>
            </section>
        </div>
        <div xmlns="http://www.w3.org/1999/xhtml" id="metrics-end"></div>
    </foreignObject>
</svg>